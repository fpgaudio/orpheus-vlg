typedef struct packed {
    integer tick_count;
} engine_state;
