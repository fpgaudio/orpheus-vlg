`default_nettype none

module mod_sum2
  ( output var signed [31:0] o_sum
  , input var signed [31:0] i_x1
  , input var signed [31:0] i_x2
  );
endmodule
